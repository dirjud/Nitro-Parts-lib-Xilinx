
`timescale  1 ps / 1 ps


module INV (O, I);

    output O;

    input  I;

	not N1 (O, I);

endmodule

