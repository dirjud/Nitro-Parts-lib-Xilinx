module BUFG (output O, input I);
   assign O=I;
endmodule

