`timescale  1 ps / 1 ps

module VCC(P);

    output P;

	assign P = 1'b1;

endmodule

