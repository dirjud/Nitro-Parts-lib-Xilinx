
`timescale  1 ps / 1 ps

module GND(G);

    output G;

	assign G = 1'b0;

endmodule

